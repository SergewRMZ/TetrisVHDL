library verilog;
use verilog.vl_types.all;
entity Tetris_vlg_vec_tst is
end Tetris_vlg_vec_tst;
