library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package Pieces_pkg is
    -- Definición de las piezas Tetris como matrices de 4x4
    type Piece_Array is array (0 to 3, 0 to 3) of std_logic;
     
    

end Pieces_pkg;
