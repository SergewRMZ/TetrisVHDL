LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE work.Pieces.ALL;
USE work.Functions.ALL;
ENTITY Tetris IS
	PORT (
		clk : IN STD_LOGIC;
		reset : IN STD_LOGIC;
		right_btn : IN STD_LOGIC;
		left_btn : IN STD_LOGIC;
		rotate_right_btn : IN STD_LOGIC;
		rotate_left_btn : IN STD_LOGIC;
		-- Salidas
		row_sel : OUT STD_LOGIC_VECTOR(0 TO 7);
		col_sel : OUT STD_LOGIC_VECTOR (0 TO 7);
		clk_desp : OUT STD_LOGIC
	);
END Tetris;

ARCHITECTURE Juego OF Tetris IS
	SIGNAL board : matrix;
	SIGNAL board_aux : matrix;

	-- State Machines
	TYPE State_Type IS (INIT, FALLING, SOLVE_COLLISION, GAME_OVER, NEXTFIGURE, ROTATION);
	SIGNAL state : State_Type := INIT;

	TYPE Action_State_Type IS (ESPERA, CLEAR, DRAW, CHARGE, DETECT_COLLISION, ROTATE_LEFT, ROTATE_RIGHT, VERIFY_LINES);
	SIGNAL state_piece : Action_State_Type := ESPERA;

	-- Matriz de Leds
	SIGNAL row_index : INTEGER := 0;

	-- Pieces
	SIGNAL current_piece : Piece_Array;
	SIGNAL next_piece : Piece_Array;

	-- Clock Signals
	SIGNAL shift_clock : STD_LOGIC := '0';
	SIGNAL init_complete : BOOLEAN := false;
	-- Seï¿½ales de debouncer
	SIGNAL right_debounced : STD_LOGIC := '0';
	SIGNAL left_debounced : STD_LOGIC := '0';
	
	SIGNAL counter_lines : INTEGER := 0;

	---------------------------------------------------------------------------------
	-- COMPONENTES
	COMPONENT Debouncer IS
		PORT (
			clk : IN STD_LOGIC;
			input_signal : IN STD_LOGIC;
			debounced_output : OUT STD_LOGIC
		);
	END COMPONENT;

	COMPONENT Divider IS
		PORT (
			clk : IN STD_LOGIC;
			clk_divider : OUT STD_LOGIC
		);
	END COMPONENT;

	---------------------------------------------------------------------------------
	-- VARIABLES COPMPARTIDAS
	SHARED VARIABLE figure_y : INTEGER RANGE 0 TO 8 := 0;
	SHARED VARIABLE figure_x : INTEGER RANGE -2 TO 8 := 0;
	---------------------------------------------------------------------------------

	---------------------------------------------------------------------------------
	----- INICIO DE LA ARQUITECTURA

BEGIN
	frecuency_divider : Divider PORT MAP(clk => clk, clk_divider => shift_clock);

	JUEGO_TETRIS : PROCESS (reset, clk, shift_clock)
		VARIABLE isCollision : BOOLEAN := false;
	BEGIN
		IF reset = '1' THEN
			REPORT "INICIANDO JUEGO";
			row_sel <= "11111111";
			FOR i IN 0 TO 7 LOOP
				FOR j IN 0 TO 7 LOOP
					board(i, j) <= '0';
					board_aux(i, j) <= '0';
				END LOOP;
			END LOOP;

			board(7, 0) <= '1';
			board(7, 1) <= '1';
			board(7, 2) <= '1';
			board(7, 3) <= '1';

			board(6, 0) <= '1';
			board(6, 1) <= '1';
			board(6, 2) <= '1';
			board(6, 3) <= '1';

			board(7, 4) <= '1';
			board(6, 4) <= '1';
			board(5, 4) <= '1';
			board(4, 4) <= '1';

			board(5, 1) <= '1';
			board(5, 2) <= '1';
			board(4, 1) <= '1';
			board(3, 1) <= '1';
			figure_x := 0;
			figure_y := 0;

			-- Cargar pieza inicial
			current_piece <= PIECE_L;

			-- Dibujar la pieza inicial en el tablero (por ejemplo, en la fila 0, columna 3)
			draw_piece(current_piece, figure_x, figure_y, board_aux);
			chargePiece(board_aux, board);

		ELSIF rising_edge(clk) THEN
		
			IF shift_clock = '1' THEN
				 figure_y := figure_y + 1;
			END IF;
			
			CASE state IS
				WHEN INIT =>
					state <= FALLING;

				WHEN FALLING =>
					CASE state_piece IS
						WHEN ESPERA =>
							state_piece <= CLEAR;

						WHEN CLEAR =>
							clearPiece(board, board_aux);
							clearMatAux(board_aux);
							state_piece <= DRAW;

						WHEN DRAW =>
							IF figure_y < 7 THEN
								draw_piece(current_piece, figure_x, figure_y, board_aux);
								state_piece <= DETECT_COLLISION;
							END IF;
						WHEN DETECT_COLLISION =>
							isCollision := check_collision(board_aux, board);
							IF NOT isCollision THEN
								state_piece <= CHARGE;

							ELSE
								REPORT "COLLISION DETECTADA" SEVERITY note;
								state <= SOLVE_COLLISION;
								state_piece <= CLEAR;
							END IF;

						WHEN CHARGE =>
							chargePiece(board_aux, board);
							REPORT "Cargando pieza en (" & INTEGER'IMAGE(figure_y) & ")" & "(" & INTEGER'IMAGE(figure_x) & ")";
							IF figure_y = 7 THEN
								state <= NEXTFIGURE;
								state_piece <= CLEAR;

							ELSE
								state_piece <= ESPERA;
							END IF;
							
						WHEN OTHERS => NULL;

					END CASE;

				WHEN NEXTFIGURE =>
					CASE state_piece IS
						WHEN CLEAR =>
							clearMatAux(board_aux);
							figure_y := 0;
							figure_x := 0;
							current_piece <= PIECE_S;
							state_piece <= DRAW;

						WHEN DRAW =>
							draw_piece(current_piece, figure_x, figure_y, board_aux);
							state_piece <= DETECT_COLLISION;
							state <= FALLING;

						WHEN OTHERS => NULL;
					END CASE;

				WHEN SOLVE_COLLISION =>
					CASE state_piece IS
						WHEN CLEAR =>
							IF figure_y > 0 THEN
								figure_y := figure_y - 1; -- Retroceder la pieza
							ELSE
								-- De estar en el estado de colision en y = 0, fin del juego.
								state <= GAME_OVER;
								REPORT "FIN DEL JUEGO";
							END IF;
							REPORT "Retrocede al ultimo estado: figure_x=" & INTEGER'IMAGE(figure_x) & ", figure_y=" & INTEGER'IMAGE(figure_y) SEVERITY note;
							clearMatAux(board_aux);
							state_piece <= DRAW;

						WHEN DRAW =>
							draw_piece(current_piece, figure_x, figure_y, board_aux);
							state_piece <= CHARGE;
 
						WHEN CHARGE =>
							chargePiece(board_aux, board);
							state_piece <= VERIFY_LINES;
							
						WHEN VERIFY_LINES => 
						   REPORT "Verificar lineas";
						   verifyLines(board, counter_lines);
						   state <= NEXTFIGURE;
							 state_piece <= CLEAR;

						WHEN OTHERS => NULL;

					END CASE;

				WHEN ROTATION =>
					CASE state_piece IS
						WHEN ROTATE_LEFT =>
							current_piece <= rotateLeft(current_piece);
							state <= FALLING;
							state_piece <= CLEAR;

						WHEN ROTATE_RIGHT =>
							current_piece <= rotateRight(current_piece);
							state <= FALLING;
							state_piece <= CLEAR;
						WHEN OTHERS => NULL;
					END CASE;

				WHEN GAME_OVER =>
					FOR i IN 0 TO 7 LOOP
						FOR j IN 0 TO 7 LOOP
							board(i, j) <= '1';
						END LOOP;
					END LOOP;
				WHEN OTHERS => NULL;
			END CASE;

			IF right_btn = '1' THEN
			   IF canMoveRight(current_piece, figure_x, figure_y, board) THEN
				    figure_x := figure_x + 1;
				  	 REPORT "Derecha -> X = " & INTEGER'IMAGE(figure_x);
			   END IF;
		  END IF;

			IF rotate_right_btn = '1' THEN
				state <= ROTATION;
				state_piece <= ROTATE_RIGHT;
			END IF;

			IF rotate_left_btn = '1' THEN
				state <= ROTATION;
			END IF;
			repaint(row_index, col_sel, row_sel, board);

		END IF;
	END PROCESS;

  PROCESS(counter_lines) IS BEGIN
    if counter_lines > 0 THEN
      REPORT "Contando lineas " & INTEGER'IMAGE(counter_lines);
    end if;
  END PROCESS; 
  
  
	clk_desp <= shift_clock;
  
END ARCHITECTURE Juego;